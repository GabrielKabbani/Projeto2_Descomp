LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

PACKAGE controls IS

  -- funct TIPO R
  CONSTANT OP_AND : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100100";
  CONSTANT OP_OR : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100101";
  CONSTANT OP_ADD : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100000";
  CONSTANT OP_SUB : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100010";
  CONSTANT OP_SLT : STD_LOGIC_VECTOR(5 DOWNTO 0) := "101010";

  constant OP_CODE_R : STD_LOGIC_VECTOR(5 downto 0) := "000000";
  -- op_code TIPO I
  CONSTANT OP_LW : STD_LOGIC_VECTOR(5 DOWNTO 0) := "100011";
  CONSTANT OP_SW : STD_LOGIC_VECTOR(5 DOWNTO 0) := "101011";
  -- op_code TIPO J
  CONSTANT OP_BEQ : STD_LOGIC_VECTOR(5 DOWNTO 0) := "000100";
  CONSTANT OP_JMP : STD_LOGIC_VECTOR(5 DOWNTO 0) := "000010";

  -- controle ULA
  CONSTANT CTRL_AND : STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
  CONSTANT CTRL_OR : STD_LOGIC_VECTOR(2 DOWNTO 0) := "001";
  CONSTANT CTRL_ADD : STD_LOGIC_VECTOR(2 DOWNTO 0) := "010";
  CONSTANT CTRL_SUB : STD_LOGIC_VECTOR(2 DOWNTO 0) := "110";
  CONSTANT CTRL_SLT : STD_LOGIC_VECTOR(2 DOWNTO 0) := "111";
--  CONSTANT CTRL_NOP : STD_LOGIC_VECTOR(2 DOWNTO 0) := "??";

  --
END PACKAGE controls;